import i2c_typedefs::*;
class random_generator extends ncsu_component;
endclass